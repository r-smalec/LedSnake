module frame_counter (

);

endmodule