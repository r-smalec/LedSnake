module prescaler_selector(
    input                   clk,
    input                   rstn,

    input                   bit_to_transmit,
    input                   all_bits_shifted,
    input                   reset_signal_finish,

    output reg              l_time_wait,
    input                   l_time_measured,
    output reg              s_time_wait,
    input                   s_time_measured,

    output reg              led_stripe_pin
);



endmodule
